** sch_path: /home/dsatizabal/simple-fet-inverter/xschem/inverter_tb.sch
**.subckt inverter_tb Vin Vout
*.ipin Vin
*.opin Vout
V1 VSS GND 1.8
X1 VSS Vin Vout VDD inverter
V2 VDD GND 0
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/sky130.lib.spice tt




Vin IN 0 pulse 0 1.8 5n 1n 1n 50n 100n
.control
tran 100p 200n
write inverter_tb.raw
.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  inverter.sym # of pins=4
** sym_path: /home/dsatizabal/simple-fet-inverter/xschem/inverter.sym
** sch_path: /home/dsatizabal/simple-fet-inverter/xschem/inverter.sch
.subckt inverter VSS IN OUT VDD
*.ipin IN
*.opin OUT
*.iopin VSS
*.iopin VDD
XM1 OUT IN VDD VDD sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VSS VSS sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
