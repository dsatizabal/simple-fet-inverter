** sch_path: /home/dsatizabal/simple-fet-inverter/xschem/custinv_tb.sch
**.subckt custinv_tb Vout
*.opin Vout
X1 net2 net1 Vout Vin custinv
V1 net1 GND 0
V2 Vin GND pulse(0 1.8 0n 1n 1n 50n 100n)
V3 net2 GND 1.8
**** begin user architecture code



.control
tran 1n 500n
write custinv_tb.raw
.endc




.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/corners/tt.spice
.include /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/dsatizabal/.volare/volare/sky130/versions/78b7bc32ddb4b6f14f76883c2e2dc5b5de9d1cbc/sky130A/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:  custinv.sym # of pins=4
** sym_path: /home/dsatizabal/simple-fet-inverter/xschem/custinv.sym
** sch_path: /home/dsatizabal/simple-fet-inverter/xschem/custinv.sch
.subckt custinv VSS VDD OUT IN
*.ipin IN
*.opin OUT
*.iopin VSS
*.iopin VDD
XM1 OUT IN VDD VDD sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT IN VSS VSS sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
